fp32log_inst : fp32log PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		result	 => result_sig
	);
