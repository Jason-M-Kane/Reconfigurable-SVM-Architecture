fp32_compare_gt_inst : fp32_compare_gt PORT MAP (
		aclr	 => aclr_sig,
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		agb	 => agb_sig
	);
