-- uart.vhd

-- Generated using ACDS version 13.0sp1 232 at 2013.11.12.05:42:32

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity uart is
	port (
		clk_clk                        : in  std_logic                     := '0';             --                        clk.clk
		reset_reset_n                  : in  std_logic                     := '0';             --                      reset.reset_n
		uart_0_external_connection_rxd : in  std_logic                     := '0';             -- uart_0_external_connection.rxd
		uart_0_external_connection_txd : out std_logic;                                        --                           .txd
		mm_bridge_0_s0_waitrequest     : out std_logic;                                        --             mm_bridge_0_s0.waitrequest
		mm_bridge_0_s0_readdata        : out std_logic_vector(31 downto 0);                    --                           .readdata
		mm_bridge_0_s0_readdatavalid   : out std_logic;                                        --                           .readdatavalid
		mm_bridge_0_s0_burstcount      : in  std_logic_vector(0 downto 0)  := (others => '0'); --                           .burstcount
		mm_bridge_0_s0_writedata       : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		mm_bridge_0_s0_address         : in  std_logic_vector(2 downto 0)  := (others => '0'); --                           .address
		mm_bridge_0_s0_write           : in  std_logic                     := '0';             --                           .write
		mm_bridge_0_s0_read            : in  std_logic                     := '0';             --                           .read
		mm_bridge_0_s0_byteenable      : in  std_logic_vector(3 downto 0)  := (others => '0'); --                           .byteenable
		mm_bridge_0_s0_debugaccess     : in  std_logic                     := '0'              --                           .debugaccess
	);
end entity uart;

architecture rtl of uart is
	component uart_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			dataavailable : out std_logic;                                        -- dataavailable
			readyfordata  : out std_logic;                                        -- readyfordata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component uart_uart_0;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			ADDRESS_WIDTH     : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(2 downto 0);                     -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_bridge;

	component altera_merlin_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(4 downto 0);                     -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_translator;

	component altera_merlin_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_chipselect            : out std_logic;                                        -- chipselect
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_translator;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	signal mm_bridge_0_m0_burstcount                                         : std_logic_vector(0 downto 0);  -- mm_bridge_0:m0_burstcount -> mm_bridge_0_m0_translator:av_burstcount
	signal mm_bridge_0_m0_waitrequest                                        : std_logic;                     -- mm_bridge_0_m0_translator:av_waitrequest -> mm_bridge_0:m0_waitrequest
	signal mm_bridge_0_m0_address                                            : std_logic_vector(2 downto 0);  -- mm_bridge_0:m0_address -> mm_bridge_0_m0_translator:av_address
	signal mm_bridge_0_m0_writedata                                          : std_logic_vector(31 downto 0); -- mm_bridge_0:m0_writedata -> mm_bridge_0_m0_translator:av_writedata
	signal mm_bridge_0_m0_write                                              : std_logic;                     -- mm_bridge_0:m0_write -> mm_bridge_0_m0_translator:av_write
	signal mm_bridge_0_m0_read                                               : std_logic;                     -- mm_bridge_0:m0_read -> mm_bridge_0_m0_translator:av_read
	signal mm_bridge_0_m0_readdata                                           : std_logic_vector(31 downto 0); -- mm_bridge_0_m0_translator:av_readdata -> mm_bridge_0:m0_readdata
	signal mm_bridge_0_m0_debugaccess                                        : std_logic;                     -- mm_bridge_0:m0_debugaccess -> mm_bridge_0_m0_translator:av_debugaccess
	signal mm_bridge_0_m0_byteenable                                         : std_logic_vector(3 downto 0);  -- mm_bridge_0:m0_byteenable -> mm_bridge_0_m0_translator:av_byteenable
	signal mm_bridge_0_m0_readdatavalid                                      : std_logic;                     -- mm_bridge_0_m0_translator:av_readdatavalid -> mm_bridge_0:m0_readdatavalid
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_waitrequest   : std_logic;                     -- uart_0_s1_translator:uav_waitrequest -> mm_bridge_0_m0_translator:uav_waitrequest
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_burstcount    : std_logic_vector(2 downto 0);  -- mm_bridge_0_m0_translator:uav_burstcount -> uart_0_s1_translator:uav_burstcount
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_writedata     : std_logic_vector(31 downto 0); -- mm_bridge_0_m0_translator:uav_writedata -> uart_0_s1_translator:uav_writedata
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_address       : std_logic_vector(4 downto 0);  -- mm_bridge_0_m0_translator:uav_address -> uart_0_s1_translator:uav_address
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_lock          : std_logic;                     -- mm_bridge_0_m0_translator:uav_lock -> uart_0_s1_translator:uav_lock
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_write         : std_logic;                     -- mm_bridge_0_m0_translator:uav_write -> uart_0_s1_translator:uav_write
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_read          : std_logic;                     -- mm_bridge_0_m0_translator:uav_read -> uart_0_s1_translator:uav_read
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_readdata      : std_logic_vector(31 downto 0); -- uart_0_s1_translator:uav_readdata -> mm_bridge_0_m0_translator:uav_readdata
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_debugaccess   : std_logic;                     -- mm_bridge_0_m0_translator:uav_debugaccess -> uart_0_s1_translator:uav_debugaccess
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_byteenable    : std_logic_vector(3 downto 0);  -- mm_bridge_0_m0_translator:uav_byteenable -> uart_0_s1_translator:uav_byteenable
	signal mm_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid : std_logic;                     -- uart_0_s1_translator:uav_readdatavalid -> mm_bridge_0_m0_translator:uav_readdatavalid
	signal uart_0_s1_translator_avalon_anti_slave_0_writedata                : std_logic_vector(15 downto 0); -- uart_0_s1_translator:av_writedata -> uart_0:writedata
	signal uart_0_s1_translator_avalon_anti_slave_0_address                  : std_logic_vector(2 downto 0);  -- uart_0_s1_translator:av_address -> uart_0:address
	signal uart_0_s1_translator_avalon_anti_slave_0_chipselect               : std_logic;                     -- uart_0_s1_translator:av_chipselect -> uart_0:chipselect
	signal uart_0_s1_translator_avalon_anti_slave_0_write                    : std_logic;                     -- uart_0_s1_translator:av_write -> uart_0_s1_translator_avalon_anti_slave_0_write:in
	signal uart_0_s1_translator_avalon_anti_slave_0_read                     : std_logic;                     -- uart_0_s1_translator:av_read -> uart_0_s1_translator_avalon_anti_slave_0_read:in
	signal uart_0_s1_translator_avalon_anti_slave_0_readdata                 : std_logic_vector(15 downto 0); -- uart_0:readdata -> uart_0_s1_translator:av_readdata
	signal uart_0_s1_translator_avalon_anti_slave_0_begintransfer            : std_logic;                     -- uart_0_s1_translator:av_begintransfer -> uart_0:begintransfer
	signal rst_controller_reset_out_reset                                    : std_logic;                     -- rst_controller:reset_out -> [mm_bridge_0:reset, mm_bridge_0_m0_translator:reset, rst_controller_reset_out_reset:in, uart_0_s1_translator:reset]
	signal reset_reset_n_ports_inv                                           : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal uart_0_s1_translator_avalon_anti_slave_0_write_ports_inv          : std_logic;                     -- uart_0_s1_translator_avalon_anti_slave_0_write:inv -> uart_0:write_n
	signal uart_0_s1_translator_avalon_anti_slave_0_read_ports_inv           : std_logic;                     -- uart_0_s1_translator_avalon_anti_slave_0_read:inv -> uart_0:read_n
	signal rst_controller_reset_out_reset_ports_inv                          : std_logic;                     -- rst_controller_reset_out_reset:inv -> uart_0:reset_n

begin

	uart_0 : component uart_uart_0
		port map (
			clk           => clk_clk,                                                  --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                 --               reset.reset_n
			address       => uart_0_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			begintransfer => uart_0_s1_translator_avalon_anti_slave_0_begintransfer,   --                    .begintransfer
			chipselect    => uart_0_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			read_n        => uart_0_s1_translator_avalon_anti_slave_0_read_ports_inv,  --                    .read_n
			write_n       => uart_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata     => uart_0_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			readdata      => uart_0_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			dataavailable => open,                                                     --                    .dataavailable
			readyfordata  => open,                                                     --                    .readyfordata
			rxd           => uart_0_external_connection_rxd,                           -- external_connection.export
			txd           => uart_0_external_connection_txd,                           --                    .export
			irq           => open                                                      --                 irq.irq
		);

	mm_bridge_0 : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			ADDRESS_WIDTH     => 3,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => clk_clk,                        --   clk.clk
			reset            => rst_controller_reset_out_reset, -- reset.reset
			s0_waitrequest   => mm_bridge_0_s0_waitrequest,     --    s0.waitrequest
			s0_readdata      => mm_bridge_0_s0_readdata,        --      .readdata
			s0_readdatavalid => mm_bridge_0_s0_readdatavalid,   --      .readdatavalid
			s0_burstcount    => mm_bridge_0_s0_burstcount,      --      .burstcount
			s0_writedata     => mm_bridge_0_s0_writedata,       --      .writedata
			s0_address       => mm_bridge_0_s0_address,         --      .address
			s0_write         => mm_bridge_0_s0_write,           --      .write
			s0_read          => mm_bridge_0_s0_read,            --      .read
			s0_byteenable    => mm_bridge_0_s0_byteenable,      --      .byteenable
			s0_debugaccess   => mm_bridge_0_s0_debugaccess,     --      .debugaccess
			m0_waitrequest   => mm_bridge_0_m0_waitrequest,     --    m0.waitrequest
			m0_readdata      => mm_bridge_0_m0_readdata,        --      .readdata
			m0_readdatavalid => mm_bridge_0_m0_readdatavalid,   --      .readdatavalid
			m0_burstcount    => mm_bridge_0_m0_burstcount,      --      .burstcount
			m0_writedata     => mm_bridge_0_m0_writedata,       --      .writedata
			m0_address       => mm_bridge_0_m0_address,         --      .address
			m0_write         => mm_bridge_0_m0_write,           --      .write
			m0_read          => mm_bridge_0_m0_read,            --      .read
			m0_byteenable    => mm_bridge_0_m0_byteenable,      --      .byteenable
			m0_debugaccess   => mm_bridge_0_m0_debugaccess      --      .debugaccess
		);

	mm_bridge_0_m0_translator : component altera_merlin_master_translator
		generic map (
			AV_ADDRESS_W                => 3,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 5,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 0,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                           --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --                     reset.reset
			uav_address              => mm_bridge_0_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => mm_bridge_0_m0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => mm_bridge_0_m0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => mm_bridge_0_m0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => mm_bridge_0_m0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => mm_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => mm_bridge_0_m0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => mm_bridge_0_m0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => mm_bridge_0_m0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => mm_bridge_0_m0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => mm_bridge_0_m0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => mm_bridge_0_m0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => mm_bridge_0_m0_waitrequest,                                        --                          .waitrequest
			av_burstcount            => mm_bridge_0_m0_burstcount,                                         --                          .burstcount
			av_byteenable            => mm_bridge_0_m0_byteenable,                                         --                          .byteenable
			av_read                  => mm_bridge_0_m0_read,                                               --                          .read
			av_readdata              => mm_bridge_0_m0_readdata,                                           --                          .readdata
			av_readdatavalid         => mm_bridge_0_m0_readdatavalid,                                      --                          .readdatavalid
			av_write                 => mm_bridge_0_m0_write,                                              --                          .write
			av_writedata             => mm_bridge_0_m0_writedata,                                          --                          .writedata
			av_debugaccess           => mm_bridge_0_m0_debugaccess,                                        --                          .debugaccess
			av_beginbursttransfer    => '0',                                                               --               (terminated)
			av_begintransfer         => '0',                                                               --               (terminated)
			av_chipselect            => '0',                                                               --               (terminated)
			av_lock                  => '0',                                                               --               (terminated)
			uav_clken                => open,                                                              --               (terminated)
			av_clken                 => '1',                                                               --               (terminated)
			uav_response             => "00",                                                              --               (terminated)
			av_response              => open,                                                              --               (terminated)
			uav_writeresponserequest => open,                                                              --               (terminated)
			uav_writeresponsevalid   => '0',                                                               --               (terminated)
			av_writeresponserequest  => '0',                                                               --               (terminated)
			av_writeresponsevalid    => open                                                               --               (terminated)
		);

	uart_0_s1_translator : component altera_merlin_slave_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 5,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                    --                    reset.reset
			uav_address              => mm_bridge_0_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => mm_bridge_0_m0_translator_avalon_universal_master_0_burstcount,    --                         .burstcount
			uav_read                 => mm_bridge_0_m0_translator_avalon_universal_master_0_read,          --                         .read
			uav_write                => mm_bridge_0_m0_translator_avalon_universal_master_0_write,         --                         .write
			uav_waitrequest          => mm_bridge_0_m0_translator_avalon_universal_master_0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => mm_bridge_0_m0_translator_avalon_universal_master_0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => mm_bridge_0_m0_translator_avalon_universal_master_0_byteenable,    --                         .byteenable
			uav_readdata             => mm_bridge_0_m0_translator_avalon_universal_master_0_readdata,      --                         .readdata
			uav_writedata            => mm_bridge_0_m0_translator_avalon_universal_master_0_writedata,     --                         .writedata
			uav_lock                 => mm_bridge_0_m0_translator_avalon_universal_master_0_lock,          --                         .lock
			uav_debugaccess          => mm_bridge_0_m0_translator_avalon_universal_master_0_debugaccess,   --                         .debugaccess
			av_address               => uart_0_s1_translator_avalon_anti_slave_0_address,                  --      avalon_anti_slave_0.address
			av_write                 => uart_0_s1_translator_avalon_anti_slave_0_write,                    --                         .write
			av_read                  => uart_0_s1_translator_avalon_anti_slave_0_read,                     --                         .read
			av_readdata              => uart_0_s1_translator_avalon_anti_slave_0_readdata,                 --                         .readdata
			av_writedata             => uart_0_s1_translator_avalon_anti_slave_0_writedata,                --                         .writedata
			av_begintransfer         => uart_0_s1_translator_avalon_anti_slave_0_begintransfer,            --                         .begintransfer
			av_chipselect            => uart_0_s1_translator_avalon_anti_slave_0_chipselect,               --                         .chipselect
			av_beginbursttransfer    => open,                                                              --              (terminated)
			av_burstcount            => open,                                                              --              (terminated)
			av_byteenable            => open,                                                              --              (terminated)
			av_readdatavalid         => '0',                                                               --              (terminated)
			av_waitrequest           => '0',                                                               --              (terminated)
			av_writebyteenable       => open,                                                              --              (terminated)
			av_lock                  => open,                                                              --              (terminated)
			av_clken                 => open,                                                              --              (terminated)
			uav_clken                => '0',                                                               --              (terminated)
			av_debugaccess           => open,                                                              --              (terminated)
			av_outputenable          => open,                                                              --              (terminated)
			uav_response             => open,                                                              --              (terminated)
			av_response              => "00",                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                              --              (terminated)
			av_writeresponserequest  => open,                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                --              (terminated)
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	uart_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not uart_0_s1_translator_avalon_anti_slave_0_write;

	uart_0_s1_translator_avalon_anti_slave_0_read_ports_inv <= not uart_0_s1_translator_avalon_anti_slave_0_read;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of uart
